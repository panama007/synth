
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity FIR is
    Port ( input    : in  STD_LOGIC;
           taps     : in  
           integer_vector;
           output   : out  STD_LOGIC);
end FIR;

architecture Behavioral of FIR is

begin


end Behavioral;

