library IEEE;
use IEEE.STD_LOGIC_1164.all;

package fonts is
    type letter is array(0 to 15) of std_logic_vector(0 to 15);
    type font_type is array(0 to 95) of letter;
    
    constant PressStart2P : font_type := (("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000111111000000","0000111111000000","0000111111000000","0000111111000000","0000111111000000","0000111111000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000000000000000","0000000000000000","0000111100000000","0000111100000000","0000000000000000","0000000000000000"),("0011110011110000","0011110011110000","0011110011110000","0011110011110000","0011110011110000","0011110011110000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0001111001111000","0001111001111000","0111111111111110","0111111111111110","0001111001111000","0001111001111000","0001111001111000","0001111001111000","0001111001111000","0001111001111000","0111111111111110","0111111111111110","0001111001111000","0001111001111000","0000000000000000","0000000000000000"),("0000000110000000","0000000110000000","0001111111111000","0001111111111000","0111100110000000","0111100110000000","0001111111111000","0001111111111000","0000000110011110","0000000110011110","0111111111111000","0111111111111000","0000000110000000","0000000110000000","0000000000000000","0000000000000000"),("0001111000000110","0001111000000110","0110011000011000","0110011000011000","0111100001100000","0111100001100000","0000000110000000","0000000110000000","0000011000011110","0000011000011110","0001100001100110","0001100001100110","0110000001111000","0110000001111000","0000000000000000","0000000000000000"),("0001111110000000","0001111110000000","0111100111100000","0111100111100000","0111100111100000","0111100111100000","0001111110000000","0001111110000000","0111100111100110","0111100111100110","0111100001111000","0111100001111000","0001111111111110","0001111111111110","0000000000000000","0000000000000000"),("0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000011110000","0000000011110000","0000001111000000","0000001111000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000001111000000","0000001111000000","0000000011110000","0000000011110000","0000000000000000","0000000000000000"),("0011110000000000","0011110000000000","0000111100000000","0000111100000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000111100000000","0000111100000000","0011110000000000","0011110000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0001111001111000","0001111001111000","0000011111100000","0000011111100000","0111111111111110","0111111111111110","0000011111100000","0000011111100000","0001111001111000","0001111001111000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0011111111111100","0011111111111100","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0011110000000000","0011110000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0011111111111100","0011111111111100","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000000000000000","0000000000000000"),("0000000000000110","0000000000000110","0000000000011000","0000000000011000","0000000001100000","0000000001100000","0000000110000000","0000000110000000","0000011000000000","0000011000000000","0001100000000000","0001100000000000","0110000000000000","0110000000000000","0000000000000000","0000000000000000"),("0000011111100000","0000011111100000","0001100001111000","0001100001111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111000011000","0001111000011000","0000011111100000","0000011111100000","0000000000000000","0000000000000000"),("0000001111000000","0000001111000000","0000111111000000","0000111111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0011111111111100","0011111111111100","0000000000000000","0000000000000000"),("0001111111111000","0001111111111000","0111100000011110","0111100000011110","0000000001111110","0000000001111110","0000011111111000","0000011111111000","0001111111100000","0001111111100000","0111111000000000","0111111000000000","0111111111111110","0111111111111110","0000000000000000","0000000000000000"),("0001111111111110","0001111111111110","0000000001111000","0000000001111000","0000000111100000","0000000111100000","0000011111111000","0000011111111000","0000000000011110","0000000000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0000000111111000","0000000111111000","0000011111111000","0000011111111000","0001111001111000","0001111001111000","0111100001111000","0111100001111000","0111111111111110","0111111111111110","0000000001111000","0000000001111000","0000000001111000","0000000001111000","0000000000000000","0000000000000000"),("0111111111111000","0111111111111000","0111100000000000","0111100000000000","0111111111111000","0111111111111000","0000000000011110","0000000000011110","0000000000011110","0000000000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0000011111111000","0000011111111000","0001111000000000","0001111000000000","0111100000000000","0111100000000000","0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0111111111111110","0111111111111110","0111100000011110","0111100000011110","0000000001111000","0000000001111000","0000000111100000","0000000111100000","0000011110000000","0000011110000000","0000011110000000","0000011110000000","0000011110000000","0000011110000000","0000000000000000","0000000000000000"),("0001111111100000","0001111111100000","0111100000011000","0111100000011000","0111111000011000","0111111000011000","0001111111100000","0001111111100000","0110000111111110","0110000111111110","0110000000011110","0110000000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0001111111111000","0001111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111110","0001111111111110","0000000000011110","0000000000011110","0000000001111000","0000000001111000","0001111111100000","0001111111100000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000000000000000","0000000000000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000000000000000","0000000000000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0011110000000000","0011110000000000","0000000000000000","0000000000000000"),("0000000011110000","0000000011110000","0000001111000000","0000001111000000","0000111100000000","0000111100000000","0011110000000000","0011110000000000","0000111100000000","0000111100000000","0000001111000000","0000001111000000","0000000011110000","0000000011110000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111111111111110","0111111111111110","0000000000000000","0000000000000000","0111111111111110","0111111111111110","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0011110000000000","0011110000000000","0000111100000000","0000111100000000","0000001111000000","0000001111000000","0000000011110000","0000000011110000","0000001111000000","0000001111000000","0000111100000000","0000111100000000","0011110000000000","0011110000000000","0000000000000000","0000000000000000"),("0001111111111000","0001111111111000","0111111111111110","0111111111111110","0111100000011110","0111100000011110","0000000001111000","0000000001111000","0000011111100000","0000011111100000","0000000000000000","0000000000000000","0000011111100000","0000011111100000","0000000000000000","0000000000000000"),("0001111111111000","0001111111111000","0110000000000110","0110000000000110","0110011111100110","0110011111100110","0110011001100110","0110011001100110","0110011111111110","0110011111111110","0110000000000000","0110000000000000","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0000011111100000","0000011111100000","0001111001111000","0001111001111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111111111111110","0111111111111110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111111111111000","0111111111111000","0000000000000000","0000000000000000"),("0000011111111000","0000011111111000","0001111000011110","0001111000011110","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0001111000011110","0001111000011110","0000011111111000","0000011111111000","0000000000000000","0000000000000000"),("0111111111100000","0111111111100000","0111100001111000","0111100001111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100001111000","0111100001111000","0111111111100000","0111111111100000","0000000000000000","0000000000000000"),("0111111111111110","0111111111111110","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111111111111000","0111111111111000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111111111111110","0111111111111110","0000000000000000","0000000000000000"),("0111111111111110","0111111111111110","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111111111111000","0111111111111000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0000000000000000","0000000000000000"),("0000011111111110","0000011111111110","0001111000000000","0001111000000000","0111100000000000","0111100000000000","0111100001111110","0111100001111110","0111100000011110","0111100000011110","0001111000011110","0001111000011110","0000011111111110","0000011111111110","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111111111111110","0111111111111110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0011111111111100","0011111111111100","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0011111111111100","0011111111111100","0000000000000000","0000000000000000"),("0000000000011110","0000000000011110","0000000000011110","0000000000011110","0000000000011110","0000000000011110","0000000000011110","0000000000011110","0000000000011110","0000000000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111100001111000","0111100001111000","0111100111100000","0111100111100000","0111111110000000","0111111110000000","0111111111100000","0111111111100000","0111100111111000","0111100111111000","0111100001111110","0111100001111110","0000000000000000","0000000000000000"),("0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011111111111100","0011111111111100","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111111001111110","0111111001111110","0111111111111110","0111111111111110","0111111111111110","0111111111111110","0111100110011110","0111100110011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111111000011110","0111111000011110","0111111110011110","0111111110011110","0111111111111110","0111111111111110","0111100111111110","0111100111111110","0111100001111110","0111100001111110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0001111111111000","0001111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111111111111000","0111111111111000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0000000000000000","0000000000000000"),("0001111111111000","0001111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100111111110","0111100111111110","0111100001111000","0111100001111000","0001111111100110","0001111111100110","0000000000000000","0000000000000000"),("0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100001111110","0111100001111110","0111111111100000","0111111111100000","0111100111111000","0111100111111000","0111100001111110","0111100001111110","0000000000000000","0000000000000000"),("0001111111100000","0001111111100000","0111100001111000","0111100001111000","0111100000000000","0111100000000000","0001111111111000","0001111111111000","0000000000011110","0000000000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0011111111111100","0011111111111100","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111111001111110","0111111001111110","0001111111111000","0001111111111000","0000011111100000","0000011111100000","0000000110000000","0000000110000000","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100110011110","0111100110011110","0111111111111110","0111111111111110","0111111111111110","0111111111111110","0111111001111110","0111111001111110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0111100000011110","0111100000011110","0111111001111110","0111111001111110","0001111111111000","0001111111111000","0000011111100000","0000011111100000","0001111111111000","0001111111111000","0111111001111110","0111111001111110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0011110000111100","0011110000111100","0011110000111100","0011110000111100","0011110000111100","0011110000111100","0000111111110000","0000111111110000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000000000000000","0000000000000000"),("0111111111111110","0111111111111110","0000000001111110","0000000001111110","0000000111111000","0000000111111000","0000011111100000","0000011111100000","0001111110000000","0001111110000000","0111111000000000","0111111000000000","0111111111111110","0111111111111110","0000000000000000","0000000000000000"),("0000111111110000","0000111111110000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000111111110000","0000111111110000","0000000000000000","0000000000000000"),("0110000000000000","0110000000000000","0001100000000000","0001100000000000","0000011000000000","0000011000000000","0000000110000000","0000000110000000","0000000001100000","0000000001100000","0000000000011000","0000000000011000","0000000000000110","0000000000000110","0000000000000000","0000000000000000"),("0011111111000000","0011111111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0011111111000000","0011111111000000","0000000000000000","0000000000000000"),("0000111111000000","0000111111000000","0011110011110000","0011110011110000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111111111111110","0111111111111110"),("0000001100000000","0000001100000000","0000000011000000","0000000011000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111111111000","0001111111111000","0000000000011110","0000000000011110","0001111111111110","0001111111111110","0111100000011110","0111100000011110","0001111111111110","0001111111111110","0000000000000000","0000000000000000"),("0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111111111110","0001111111111110","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111100000000000","0001111111111110","0001111111111110","0000000000000000","0000000000000000"),("0000000000011110","0000000000011110","0000000000011110","0000000000011110","0001111111111110","0001111111111110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111110","0001111111111110","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111111111000","0001111111111000","0111100000011110","0111100000011110","0111111111111110","0111111111111110","0111100000000000","0111100000000000","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0000000011111100","0000000011111100","0000001111000000","0000001111000000","0011111111111100","0011111111111100","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111111111110","0001111111111110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111110","0001111111111110","0000000000011110","0000000000011110","0001111111111000","0001111111111000"),("0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0000001111000000","0000001111000000","0000000000000000","0000000000000000","0000111111000000","0000111111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0011111111111100","0011111111111100","0000000000000000","0000000000000000"),("0000000011110000","0000000011110000","0000000000000000","0000000000000000","0000001111110000","0000001111110000","0000000011110000","0000000011110000","0000000011110000","0000000011110000","0000000011110000","0000000011110000","0000000011110000","0000000011110000","0011111111000000","0011111111000000"),("0111100000000000","0111100000000000","0111100000000000","0111100000000000","0111100001111110","0111100001111110","0111111111111000","0111111111111000","0111111111100000","0111111111100000","0111100111111000","0111100111111000","0111100001111110","0111100001111110","0000000000000000","0000000000000000"),("0000111111000000","0000111111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0011111111111100","0011111111111100","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111111111111000","0111111111111000","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111111111000","0001111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111000","0001111111111000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111111111111000","0111111111111000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111111111111000","0111111111111000","0111100000000000","0111100000000000","0111100000000000","0111100000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111111111110","0001111111111110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111110","0001111111111110","0000000000011110","0000000000011110","0000000000011110","0000000000011110"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0011110011111100","0011110011111100","0011111100000000","0011111100000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0011110000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111111111000","0001111111111000","0111100000000000","0111100000000000","0001111111111000","0001111111111000","0000000000011110","0000000000011110","0111111111111000","0111111111111000","0000000000000000","0000000000000000"),("0000001111000000","0000001111000000","0000001111000000","0000001111000000","0011111111111100","0011111111111100","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111110","0001111111111110","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0011110000111100","0011110000111100","0011110000111100","0011110000111100","0011110000111100","0011110000111100","0000111111110000","0000111111110000","0000001111000000","0000001111000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0110011110011110","0001111111111110","0001111111111110","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111100000011110","0111100000011110","0111111111111110","0111111111111110","0000011111100000","0000011111100000","0111111111111110","0111111111111110","0111100000011110","0111100000011110","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0111100000011110","0001111111111110","0001111111111110","0000000000011110","0000000000011110","0001111111111000","0001111111111000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0111111111111110","0111111111111110","0000000111111000","0000000111111000","0000011111100000","0000011111100000","0001111110000000","0001111110000000","0111111111111110","0111111111111110","0000000000000000","0000000000000000"),("0000000011110000","0000000011110000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000111100000000","0000111100000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000000011110000","0000000011110000","0000000000000000","0000000000000000"),("0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000001111000000","0000000000000000","0000000000000000"),("0011110000000000","0011110000000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0000001111000000","0000001111000000","0000111100000000","0000111100000000","0000111100000000","0000111100000000","0011110000000000","0011110000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0001111110000000","0001111110000000","0110011111100110","0110011111100110","0000000111111000","0000000111111000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000"),("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0011110011110000","0011110011110000","0011110011110000","0011110011110000","0000000000000000","0000000000000000"));

    constant font : font_type := PressStart2P;
end package fonts;
