
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity parameter_controller is
--    generic ( pages : integer := 2;
--              controls: integer := 4);
--    port ( clk     : in std_logic;
--           rotaries_in: in rotaries_array(0 to controls);
--           speaker : out std_logic;
--           cathodes: out std_logic_vector(6 downto 0);
--           anodes  : inout std_logic_vector(3 downto 0));
end parameter_controller;

architecture Behavioral of parameter_controller is

begin


end Behavioral;

